module pipeline
#()
(

);


endmodule
